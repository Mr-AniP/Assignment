module vdf_3_a(CLK, A, B, C, D, E, OUT);
input CLK;
input A;
input B;
input C;
input D;
input E;
output OUT;
wire CLK;
wire A;
wire B;
wire C;
wire D;
wire E;
wire OUT;
wire _0000_;
wire _0001_;
wire _0010_;
wire _0011_;
wire _0100_;
wire _0101_;
wire _0110_;
wire _0111_;
wire _1000_;
NAND2_X1 N1(.A1(D),.A2(E),.ZN(_0000_));
DFF_X1 F1(.D(_0000_),.CK(CLK),.Q(_0001_),.QN(_0010_));
AND2_X1 A1(.A1(C),.A2(_0001_),.ZN(_0011_));
DFF_X1 F2(.D(_0011_),.CK(CLK),.Q(_0100_),.QN(_0101_));
AND2_X1 A2(.A1(B),.A2(_0100_),.ZN(_0110_));
DFF_X1 F3(.D(_0110_),.CK(CLK),.Q(_0111_),.QN(_1000_));
AND2_X1 A3(.A1(A),.A2(_0111_),.ZN(Q));
endmodule