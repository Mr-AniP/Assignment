module vdf_3_b(CLK, A, B, C, D, E, SI, SE, OUT, SO);
input CLK;
input A;
input B;
input C;
input D;
input E;
input SI;
input SE;
output OUT;
output SO;
wire CLK;
wire A;
wire B;
wire C;
wire D;
wire E;
wire SI;
wire SE;
wire OUT;
wire SO;
wire _000_;
wire _001_;
wire _010_;
wire _011_;
wire _100_;
wire _101_;
wire _110_;
wire _111_;
NAND2_X1 N1(.A1(D),.A2(E),.ZN(_000_));
SDFF_X1 F1(.D(_000_),.SE(SE),.SI(SI),.CK(CLK),.Q(_001_),.QN(_010_));
AND2_X1 A1(.A1(C),.A2(_001_),.ZN(_011_));
SDFF_X1 F2(.D(_011_),.SE(SE),.SI(_001_),.CK(CLK),.Q(_100_),.QN(_101_));
AND2_X1 A2(.A1(B),.A2(_100_),.ZN(_110_));
SDFF_X1 F3(.D(_110_),.SE(SE),.SI(_100_),.CK(CLK),.Q(SO),.QN(_111_));
AND2_X1 A3(.A1(A),.A2(SO),.ZN(Q));
endmodule